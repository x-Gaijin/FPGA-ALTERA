module division(
input [2:0]a,
input[2:0]b,
output[2:0]division
);
assign division = a/b;
endmodule
