module multiplication(
input [2:0]a,
input[2:0]b,
output[4:0]multiply
);
assign multiply = a*b;
endmodule
