module notequal(
input [2:0]a,
input[2:0]b,
output result
);
assign result = (a!=b);
endmodule
