module subtraction(
input [2:0]a,
input [2:0]b,
output [2:0]subtract

);

assign subtract = a-b;
endmodule